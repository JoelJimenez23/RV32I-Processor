module controller();



endmodule
